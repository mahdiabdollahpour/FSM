library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
   entity sine_cosine is
       generic(M: natural :=32);
   Port(
	clk : in std_logic;
	reset : in std_logic;
   degree: in std_logic_vector(11 downto 0);
   sine: out std_logic_vector(M - 1 downto 0);
   cosine: out std_logic_vector(M - 1 downto 0)
);
   end sine_cosine;
   architecture Behavioral of sine_cosine is
   
       signal cout : std_logic;
   begin
   
       process(degree, clk)
       begin
		 if(falling_edge(clk)) then
       case degree is
       when X"000" => cosine <= X"00001000";
       when X"001" => cosine <= X"00000FFF";
       when X"002" => cosine <= X"00000FFD";
       when X"003" => cosine <= X"00000FFA";
       when X"004" => cosine <= X"00000FF6";
       when X"005" => cosine <= X"00000FF0";
       when X"006" => cosine <= X"00000FE9";
       when X"007" => cosine <= X"00000FE1";
       when X"008" => cosine <= X"00000FD8";
       when X"009" => cosine <= X"00000FCD";
       when X"00A" => cosine <= X"00000FC1";
       when X"00B" => cosine <= X"00000FB4";
       when X"00C" => cosine <= X"00000FA6";
       when X"00D" => cosine <= X"00000F97";
       when X"00E" => cosine <= X"00000F86";
       when X"00F" => cosine <= X"00000F74";
       when X"010" => cosine <= X"00000F61";
       when X"011" => cosine <= X"00000F4D";
       when X"012" => cosine <= X"00000F37";
       when X"013" => cosine <= X"00000F20";
       when X"014" => cosine <= X"00000F08";
       when X"015" => cosine <= X"00000EEF";
       when X"016" => cosine <= X"00000ED5";
       when X"017" => cosine <= X"00000EBA";
       when X"018" => cosine <= X"00000E9D";
       when X"019" => cosine <= X"00000E80";
       when X"01A" => cosine <= X"00000E61";
       when X"01B" => cosine <= X"00000E41";
       when X"01C" => cosine <= X"00000E20";
       when X"01D" => cosine <= X"00000DFE";
       when X"01E" => cosine <= X"00000DDB";
       when X"01F" => cosine <= X"00000DB6";
       when X"020" => cosine <= X"00000D91";
       when X"021" => cosine <= X"00000D6B";
       when X"022" => cosine <= X"00000D43";
       when X"023" => cosine <= X"00000D1B";
       when X"024" => cosine <= X"00000CF1";
       when X"025" => cosine <= X"00000CC7";
       when X"026" => cosine <= X"00000C9B";
       when X"027" => cosine <= X"00000C6F";
       when X"028" => cosine <= X"00000C41";
       when X"029" => cosine <= X"00000C13";
       when X"02A" => cosine <= X"00000BE3";
       when X"02B" => cosine <= X"00000BB3";
       when X"02C" => cosine <= X"00000B82";
       when X"02D" => cosine <= X"00000B50";
       when X"02E" => cosine <= X"00000B1D";
       when X"02F" => cosine <= X"00000AE9";
       when X"030" => cosine <= X"00000AB4";
       when X"031" => cosine <= X"00000A7F";
       when X"032" => cosine <= X"00000A48";
       when X"033" => cosine <= X"00000A11";
       when X"034" => cosine <= X"000009D9";
       when X"035" => cosine <= X"000009A1";
       when X"036" => cosine <= X"00000967";
       when X"037" => cosine <= X"0000092D";
       when X"038" => cosine <= X"000008F2";
       when X"039" => cosine <= X"000008B6";
       when X"03A" => cosine <= X"0000087A";
       when X"03B" => cosine <= X"0000083D";
       when X"03C" => cosine <= X"00000800";
       when X"03D" => cosine <= X"000007C1";
       when X"03E" => cosine <= X"00000782";
       when X"03F" => cosine <= X"00000743";
       when X"040" => cosine <= X"00000703";
       when X"041" => cosine <= X"000006C3";
       when X"042" => cosine <= X"00000681";
       when X"043" => cosine <= X"00000640";
       when X"044" => cosine <= X"000005FE";
       when X"045" => cosine <= X"000005BB";
       when X"046" => cosine <= X"00000578";
       when X"047" => cosine <= X"00000535";
       when X"048" => cosine <= X"000004F1";
       when X"049" => cosine <= X"000004AD";
       when X"04A" => cosine <= X"00000469";
       when X"04B" => cosine <= X"00000424";
       when X"04C" => cosine <= X"000003DE";
       when X"04D" => cosine <= X"00000399";
       when X"04E" => cosine <= X"00000353";
       when X"04F" => cosine <= X"0000030D";
       when X"050" => cosine <= X"000002C7";
       when X"051" => cosine <= X"00000280";
       when X"052" => cosine <= X"0000023A";
       when X"053" => cosine <= X"000001F3";
       when X"054" => cosine <= X"000001AC";
       when X"055" => cosine <= X"00000164";
       when X"056" => cosine <= X"0000011D";
       when X"057" => cosine <= X"000000D6";
       when X"058" => cosine <= X"0000008E";
       when X"059" => cosine <= X"00000047";
       when X"05A" => cosine <= X"00000000";
       when X"05B" => cosine <= X"FFFFFFB9";
       when X"05C" => cosine <= X"FFFFFF72";
       when X"05D" => cosine <= X"FFFFFF2A";
       when X"05E" => cosine <= X"FFFFFEE3";
       when X"05F" => cosine <= X"FFFFFE9C";
       when X"060" => cosine <= X"FFFFFE54";
       when X"061" => cosine <= X"FFFFFE0D";
       when X"062" => cosine <= X"FFFFFDC6";
       when X"063" => cosine <= X"FFFFFD80";
       when X"064" => cosine <= X"FFFFFD39";
       when X"065" => cosine <= X"FFFFFCF3";
       when X"066" => cosine <= X"FFFFFCAD";
       when X"067" => cosine <= X"FFFFFC67";
       when X"068" => cosine <= X"FFFFFC22";
       when X"069" => cosine <= X"FFFFFBDC";
       when X"06A" => cosine <= X"FFFFFB97";
       when X"06B" => cosine <= X"FFFFFB53";
       when X"06C" => cosine <= X"FFFFFB0F";
       when X"06D" => cosine <= X"FFFFFACB";
       when X"06E" => cosine <= X"FFFFFA88";
       when X"06F" => cosine <= X"FFFFFA45";
       when X"070" => cosine <= X"FFFFFA02";
       when X"071" => cosine <= X"FFFFF9C0";
       when X"072" => cosine <= X"FFFFF97F";
       when X"073" => cosine <= X"FFFFF93D";
       when X"074" => cosine <= X"FFFFF8FD";
       when X"075" => cosine <= X"FFFFF8BD";
       when X"076" => cosine <= X"FFFFF87E";
       when X"077" => cosine <= X"FFFFF83F";
       when X"078" => cosine <= X"FFFFF801";
       when X"079" => cosine <= X"FFFFF7C3";
       when X"07A" => cosine <= X"FFFFF786";
       when X"07B" => cosine <= X"FFFFF74A";
       when X"07C" => cosine <= X"FFFFF70E";
       when X"07D" => cosine <= X"FFFFF6D3";
       when X"07E" => cosine <= X"FFFFF699";
       when X"07F" => cosine <= X"FFFFF65F";
       when X"080" => cosine <= X"FFFFF627";
       when X"081" => cosine <= X"FFFFF5EF";
       when X"082" => cosine <= X"FFFFF5B8";
       when X"083" => cosine <= X"FFFFF581";
       when X"084" => cosine <= X"FFFFF54C";
       when X"085" => cosine <= X"FFFFF517";
       when X"086" => cosine <= X"FFFFF4E3";
       when X"087" => cosine <= X"FFFFF4B0";
       when X"088" => cosine <= X"FFFFF47E";
       when X"089" => cosine <= X"FFFFF44D";
       when X"08A" => cosine <= X"FFFFF41D";
       when X"08B" => cosine <= X"FFFFF3ED";
       when X"08C" => cosine <= X"FFFFF3BF";
       when X"08D" => cosine <= X"FFFFF391";
       when X"08E" => cosine <= X"FFFFF365";
       when X"08F" => cosine <= X"FFFFF339";
       when X"090" => cosine <= X"FFFFF30F";
       when X"091" => cosine <= X"FFFFF2E5";
       when X"092" => cosine <= X"FFFFF2BD";
       when X"093" => cosine <= X"FFFFF295";
       when X"094" => cosine <= X"FFFFF26F";
       when X"095" => cosine <= X"FFFFF24A";
       when X"096" => cosine <= X"FFFFF225";
       when X"097" => cosine <= X"FFFFF202";
       when X"098" => cosine <= X"FFFFF1E0";
       when X"099" => cosine <= X"FFFFF1BF";
       when X"09A" => cosine <= X"FFFFF19F";
       when X"09B" => cosine <= X"FFFFF180";
       when X"09C" => cosine <= X"FFFFF163";
       when X"09D" => cosine <= X"FFFFF146";
       when X"09E" => cosine <= X"FFFFF12B";
       when X"09F" => cosine <= X"FFFFF111";
       when X"0A0" => cosine <= X"FFFFF0F8";
       when X"0A1" => cosine <= X"FFFFF0E0";
       when X"0A2" => cosine <= X"FFFFF0C9";
       when X"0A3" => cosine <= X"FFFFF0B3";
       when X"0A4" => cosine <= X"FFFFF09F";
       when X"0A5" => cosine <= X"FFFFF08C";
       when X"0A6" => cosine <= X"FFFFF07A";
       when X"0A7" => cosine <= X"FFFFF069";
       when X"0A8" => cosine <= X"FFFFF05A";
       when X"0A9" => cosine <= X"FFFFF04C";
       when X"0AA" => cosine <= X"FFFFF03F";
       when X"0AB" => cosine <= X"FFFFF033";
       when X"0AC" => cosine <= X"FFFFF028";
       when X"0AD" => cosine <= X"FFFFF01F";
       when X"0AE" => cosine <= X"FFFFF017";
       when X"0AF" => cosine <= X"FFFFF010";
       when X"0B0" => cosine <= X"FFFFF00A";
       when X"0B1" => cosine <= X"FFFFF006";
       when X"0B2" => cosine <= X"FFFFF003";
       when X"0B3" => cosine <= X"FFFFF001";
       when X"0B4" => cosine <= X"FFFFF000";
       when X"0B5" => cosine <= X"FFFFF001";
       when X"0B6" => cosine <= X"FFFFF003";
       when X"0B7" => cosine <= X"FFFFF006";
       when X"0B8" => cosine <= X"FFFFF00A";
       when X"0B9" => cosine <= X"FFFFF010";
       when X"0BA" => cosine <= X"FFFFF017";
       when X"0BB" => cosine <= X"FFFFF01F";
       when X"0BC" => cosine <= X"FFFFF028";
       when X"0BD" => cosine <= X"FFFFF033";
       when X"0BE" => cosine <= X"FFFFF03F";
       when X"0BF" => cosine <= X"FFFFF04C";
       when X"0C0" => cosine <= X"FFFFF05A";
       when X"0C1" => cosine <= X"FFFFF069";
       when X"0C2" => cosine <= X"FFFFF07A";
       when X"0C3" => cosine <= X"FFFFF08C";
       when X"0C4" => cosine <= X"FFFFF09F";
       when X"0C5" => cosine <= X"FFFFF0B3";
       when X"0C6" => cosine <= X"FFFFF0C9";
       when X"0C7" => cosine <= X"FFFFF0E0";
       when X"0C8" => cosine <= X"FFFFF0F8";
       when X"0C9" => cosine <= X"FFFFF111";
       when X"0CA" => cosine <= X"FFFFF12B";
       when X"0CB" => cosine <= X"FFFFF146";
       when X"0CC" => cosine <= X"FFFFF163";
       when X"0CD" => cosine <= X"FFFFF180";
       when X"0CE" => cosine <= X"FFFFF19F";
       when X"0CF" => cosine <= X"FFFFF1BF";
       when X"0D0" => cosine <= X"FFFFF1E0";
       when X"0D1" => cosine <= X"FFFFF202";
       when X"0D2" => cosine <= X"FFFFF225";
       when X"0D3" => cosine <= X"FFFFF24A";
       when X"0D4" => cosine <= X"FFFFF26F";
       when X"0D5" => cosine <= X"FFFFF295";
       when X"0D6" => cosine <= X"FFFFF2BD";
       when X"0D7" => cosine <= X"FFFFF2E5";
       when X"0D8" => cosine <= X"FFFFF30F";
       when X"0D9" => cosine <= X"FFFFF339";
       when X"0DA" => cosine <= X"FFFFF365";
       when X"0DB" => cosine <= X"FFFFF391";
       when X"0DC" => cosine <= X"FFFFF3BF";
       when X"0DD" => cosine <= X"FFFFF3ED";
       when X"0DE" => cosine <= X"FFFFF41D";
       when X"0DF" => cosine <= X"FFFFF44D";
       when X"0E0" => cosine <= X"FFFFF47E";
       when X"0E1" => cosine <= X"FFFFF4B0";
       when X"0E2" => cosine <= X"FFFFF4E3";
       when X"0E3" => cosine <= X"FFFFF517";
       when X"0E4" => cosine <= X"FFFFF54C";
       when X"0E5" => cosine <= X"FFFFF581";
       when X"0E6" => cosine <= X"FFFFF5B8";
       when X"0E7" => cosine <= X"FFFFF5EF";
       when X"0E8" => cosine <= X"FFFFF627";
       when X"0E9" => cosine <= X"FFFFF65F";
       when X"0EA" => cosine <= X"FFFFF699";
       when X"0EB" => cosine <= X"FFFFF6D3";
       when X"0EC" => cosine <= X"FFFFF70E";
       when X"0ED" => cosine <= X"FFFFF74A";
       when X"0EE" => cosine <= X"FFFFF786";
       when X"0EF" => cosine <= X"FFFFF7C3";
       when X"0F0" => cosine <= X"FFFFF800";
       when X"0F1" => cosine <= X"FFFFF83F";
       when X"0F2" => cosine <= X"FFFFF87E";
       when X"0F3" => cosine <= X"FFFFF8BD";
       when X"0F4" => cosine <= X"FFFFF8FD";
       when X"0F5" => cosine <= X"FFFFF93D";
       when X"0F6" => cosine <= X"FFFFF97F";
       when X"0F7" => cosine <= X"FFFFF9C0";
       when X"0F8" => cosine <= X"FFFFFA02";
       when X"0F9" => cosine <= X"FFFFFA45";
       when X"0FA" => cosine <= X"FFFFFA88";
       when X"0FB" => cosine <= X"FFFFFACB";
       when X"0FC" => cosine <= X"FFFFFB0F";
       when X"0FD" => cosine <= X"FFFFFB53";
       when X"0FE" => cosine <= X"FFFFFB97";
       when X"0FF" => cosine <= X"FFFFFBDC";
       when X"100" => cosine <= X"FFFFFC22";
       when X"101" => cosine <= X"FFFFFC67";
       when X"102" => cosine <= X"FFFFFCAD";
       when X"103" => cosine <= X"FFFFFCF3";
       when X"104" => cosine <= X"FFFFFD39";
       when X"105" => cosine <= X"FFFFFD80";
       when X"106" => cosine <= X"FFFFFDC6";
       when X"107" => cosine <= X"FFFFFE0D";
       when X"108" => cosine <= X"FFFFFE54";
       when X"109" => cosine <= X"FFFFFE9C";
       when X"10A" => cosine <= X"FFFFFEE3";
       when X"10B" => cosine <= X"FFFFFF2A";
       when X"10C" => cosine <= X"FFFFFF72";
       when X"10D" => cosine <= X"FFFFFFB9";
       when X"10E" => cosine <= X"00000000";
       when X"10F" => cosine <= X"00000047";
       when X"110" => cosine <= X"0000008E";
       when X"111" => cosine <= X"000000D6";
       when X"112" => cosine <= X"0000011D";
       when X"113" => cosine <= X"00000164";
       when X"114" => cosine <= X"000001AC";
       when X"115" => cosine <= X"000001F3";
       when X"116" => cosine <= X"0000023A";
       when X"117" => cosine <= X"00000280";
       when X"118" => cosine <= X"000002C7";
       when X"119" => cosine <= X"0000030D";
       when X"11A" => cosine <= X"00000353";
       when X"11B" => cosine <= X"00000399";
       when X"11C" => cosine <= X"000003DE";
       when X"11D" => cosine <= X"00000424";
       when X"11E" => cosine <= X"00000469";
       when X"11F" => cosine <= X"000004AD";
       when X"120" => cosine <= X"000004F1";
       when X"121" => cosine <= X"00000535";
       when X"122" => cosine <= X"00000578";
       when X"123" => cosine <= X"000005BB";
       when X"124" => cosine <= X"000005FE";
       when X"125" => cosine <= X"00000640";
       when X"126" => cosine <= X"00000681";
       when X"127" => cosine <= X"000006C3";
       when X"128" => cosine <= X"00000703";
       when X"129" => cosine <= X"00000743";
       when X"12A" => cosine <= X"00000782";
       when X"12B" => cosine <= X"000007C1";
       when X"12C" => cosine <= X"00000800";
       when X"12D" => cosine <= X"0000083D";
       when X"12E" => cosine <= X"0000087A";
       when X"12F" => cosine <= X"000008B6";
       when X"130" => cosine <= X"000008F2";
       when X"131" => cosine <= X"0000092D";
       when X"132" => cosine <= X"00000967";
       when X"133" => cosine <= X"000009A1";
       when X"134" => cosine <= X"000009D9";
       when X"135" => cosine <= X"00000A11";
       when X"136" => cosine <= X"00000A48";
       when X"137" => cosine <= X"00000A7F";
       when X"138" => cosine <= X"00000AB4";
       when X"139" => cosine <= X"00000AE9";
       when X"13A" => cosine <= X"00000B1D";
       when X"13B" => cosine <= X"00000B50";
       when X"13C" => cosine <= X"00000B82";
       when X"13D" => cosine <= X"00000BB3";
       when X"13E" => cosine <= X"00000BE3";
       when X"13F" => cosine <= X"00000C13";
       when X"140" => cosine <= X"00000C41";
       when X"141" => cosine <= X"00000C6F";
       when X"142" => cosine <= X"00000C9B";
       when X"143" => cosine <= X"00000CC7";
       when X"144" => cosine <= X"00000CF1";
       when X"145" => cosine <= X"00000D1B";
       when X"146" => cosine <= X"00000D43";
       when X"147" => cosine <= X"00000D6B";
       when X"148" => cosine <= X"00000D91";
       when X"149" => cosine <= X"00000DB6";
       when X"14A" => cosine <= X"00000DDB";
       when X"14B" => cosine <= X"00000DFE";
       when X"14C" => cosine <= X"00000E20";
       when X"14D" => cosine <= X"00000E41";
       when X"14E" => cosine <= X"00000E61";
       when X"14F" => cosine <= X"00000E80";
       when X"150" => cosine <= X"00000E9D";
       when X"151" => cosine <= X"00000EBA";
       when X"152" => cosine <= X"00000ED5";
       when X"153" => cosine <= X"00000EEF";
       when X"154" => cosine <= X"00000F08";
       when X"155" => cosine <= X"00000F20";
       when X"156" => cosine <= X"00000F37";
       when X"157" => cosine <= X"00000F4D";
       when X"158" => cosine <= X"00000F61";
       when X"159" => cosine <= X"00000F74";
       when X"15A" => cosine <= X"00000F86";
       when X"15B" => cosine <= X"00000F97";
       when X"15C" => cosine <= X"00000FA6";
       when X"15D" => cosine <= X"00000FB4";
       when X"15E" => cosine <= X"00000FC1";
       when X"15F" => cosine <= X"00000FCD";
       when X"160" => cosine <= X"00000FD8";
       when X"161" => cosine <= X"00000FE1";
       when X"162" => cosine <= X"00000FE9";
       when X"163" => cosine <= X"00000FF0";
       when X"164" => cosine <= X"00000FF6";
       when X"165" => cosine <= X"00000FFA";
       when X"166" => cosine <= X"00000FFD";
       when X"167" => cosine <= X"00000FFF";
       when X"168" => cosine <= X"00001000";
       when others => cosine <= X"FFFFFFFF";
       end case;
       case degree is
       when X"000" => sine <= X"00000000";
       when X"001" => sine <= X"00000047";
       when X"002" => sine <= X"0000008E";
       when X"003" => sine <= X"000000D6";
       when X"004" => sine <= X"0000011D";
       when X"005" => sine <= X"00000164";
       when X"006" => sine <= X"000001AC";
       when X"007" => sine <= X"000001F3";
       when X"008" => sine <= X"0000023A";
       when X"009" => sine <= X"00000280";
       when X"00A" => sine <= X"000002C7";
       when X"00B" => sine <= X"0000030D";
       when X"00C" => sine <= X"00000353";
       when X"00D" => sine <= X"00000399";
       when X"00E" => sine <= X"000003DE";
       when X"00F" => sine <= X"00000424";
       when X"010" => sine <= X"00000469";
       when X"011" => sine <= X"000004AD";
       when X"012" => sine <= X"000004F1";
       when X"013" => sine <= X"00000535";
       when X"014" => sine <= X"00000578";
       when X"015" => sine <= X"000005BB";
       when X"016" => sine <= X"000005FE";
       when X"017" => sine <= X"00000640";
       when X"018" => sine <= X"00000681";
       when X"019" => sine <= X"000006C3";
       when X"01A" => sine <= X"00000703";
       when X"01B" => sine <= X"00000743";
       when X"01C" => sine <= X"00000782";
       when X"01D" => sine <= X"000007C1";
       when X"01E" => sine <= X"000007FF";
       when X"01F" => sine <= X"0000083D";
       when X"020" => sine <= X"0000087A";
       when X"021" => sine <= X"000008B6";
       when X"022" => sine <= X"000008F2";
       when X"023" => sine <= X"0000092D";
       when X"024" => sine <= X"00000967";
       when X"025" => sine <= X"000009A1";
       when X"026" => sine <= X"000009D9";
       when X"027" => sine <= X"00000A11";
       when X"028" => sine <= X"00000A48";
       when X"029" => sine <= X"00000A7F";
       when X"02A" => sine <= X"00000AB4";
       when X"02B" => sine <= X"00000AE9";
       when X"02C" => sine <= X"00000B1D";
       when X"02D" => sine <= X"00000B50";
       when X"02E" => sine <= X"00000B82";
       when X"02F" => sine <= X"00000BB3";
       when X"030" => sine <= X"00000BE3";
       when X"031" => sine <= X"00000C13";
       when X"032" => sine <= X"00000C41";
       when X"033" => sine <= X"00000C6F";
       when X"034" => sine <= X"00000C9B";
       when X"035" => sine <= X"00000CC7";
       when X"036" => sine <= X"00000CF1";
       when X"037" => sine <= X"00000D1B";
       when X"038" => sine <= X"00000D43";
       when X"039" => sine <= X"00000D6B";
       when X"03A" => sine <= X"00000D91";
       when X"03B" => sine <= X"00000DB6";
       when X"03C" => sine <= X"00000DDB";
       when X"03D" => sine <= X"00000DFE";
       when X"03E" => sine <= X"00000E20";
       when X"03F" => sine <= X"00000E41";
       when X"040" => sine <= X"00000E61";
       when X"041" => sine <= X"00000E80";
       when X"042" => sine <= X"00000E9D";
       when X"043" => sine <= X"00000EBA";
       when X"044" => sine <= X"00000ED5";
       when X"045" => sine <= X"00000EEF";
       when X"046" => sine <= X"00000F08";
       when X"047" => sine <= X"00000F20";
       when X"048" => sine <= X"00000F37";
       when X"049" => sine <= X"00000F4D";
       when X"04A" => sine <= X"00000F61";
       when X"04B" => sine <= X"00000F74";
       when X"04C" => sine <= X"00000F86";
       when X"04D" => sine <= X"00000F97";
       when X"04E" => sine <= X"00000FA6";
       when X"04F" => sine <= X"00000FB4";
       when X"050" => sine <= X"00000FC1";
       when X"051" => sine <= X"00000FCD";
       when X"052" => sine <= X"00000FD8";
       when X"053" => sine <= X"00000FE1";
       when X"054" => sine <= X"00000FE9";
       when X"055" => sine <= X"00000FF0";
       when X"056" => sine <= X"00000FF6";
       when X"057" => sine <= X"00000FFA";
       when X"058" => sine <= X"00000FFD";
       when X"059" => sine <= X"00000FFF";
       when X"05A" => sine <= X"00001000";
       when X"05B" => sine <= X"00000FFF";
       when X"05C" => sine <= X"00000FFD";
       when X"05D" => sine <= X"00000FFA";
       when X"05E" => sine <= X"00000FF6";
       when X"05F" => sine <= X"00000FF0";
       when X"060" => sine <= X"00000FE9";
       when X"061" => sine <= X"00000FE1";
       when X"062" => sine <= X"00000FD8";
       when X"063" => sine <= X"00000FCD";
       when X"064" => sine <= X"00000FC1";
       when X"065" => sine <= X"00000FB4";
       when X"066" => sine <= X"00000FA6";
       when X"067" => sine <= X"00000F97";
       when X"068" => sine <= X"00000F86";
       when X"069" => sine <= X"00000F74";
       when X"06A" => sine <= X"00000F61";
       when X"06B" => sine <= X"00000F4D";
       when X"06C" => sine <= X"00000F37";
       when X"06D" => sine <= X"00000F20";
       when X"06E" => sine <= X"00000F08";
       when X"06F" => sine <= X"00000EEF";
       when X"070" => sine <= X"00000ED5";
       when X"071" => sine <= X"00000EBA";
       when X"072" => sine <= X"00000E9D";
       when X"073" => sine <= X"00000E80";
       when X"074" => sine <= X"00000E61";
       when X"075" => sine <= X"00000E41";
       when X"076" => sine <= X"00000E20";
       when X"077" => sine <= X"00000DFE";
       when X"078" => sine <= X"00000DDB";
       when X"079" => sine <= X"00000DB6";
       when X"07A" => sine <= X"00000D91";
       when X"07B" => sine <= X"00000D6B";
       when X"07C" => sine <= X"00000D43";
       when X"07D" => sine <= X"00000D1B";
       when X"07E" => sine <= X"00000CF1";
       when X"07F" => sine <= X"00000CC7";
       when X"080" => sine <= X"00000C9B";
       when X"081" => sine <= X"00000C6F";
       when X"082" => sine <= X"00000C41";
       when X"083" => sine <= X"00000C13";
       when X"084" => sine <= X"00000BE3";
       when X"085" => sine <= X"00000BB3";
       when X"086" => sine <= X"00000B82";
       when X"087" => sine <= X"00000B50";
       when X"088" => sine <= X"00000B1D";
       when X"089" => sine <= X"00000AE9";
       when X"08A" => sine <= X"00000AB4";
       when X"08B" => sine <= X"00000A7F";
       when X"08C" => sine <= X"00000A48";
       when X"08D" => sine <= X"00000A11";
       when X"08E" => sine <= X"000009D9";
       when X"08F" => sine <= X"000009A1";
       when X"090" => sine <= X"00000967";
       when X"091" => sine <= X"0000092D";
       when X"092" => sine <= X"000008F2";
       when X"093" => sine <= X"000008B6";
       when X"094" => sine <= X"0000087A";
       when X"095" => sine <= X"0000083D";
       when X"096" => sine <= X"000007FF";
       when X"097" => sine <= X"000007C1";
       when X"098" => sine <= X"00000782";
       when X"099" => sine <= X"00000743";
       when X"09A" => sine <= X"00000703";
       when X"09B" => sine <= X"000006C3";
       when X"09C" => sine <= X"00000681";
       when X"09D" => sine <= X"00000640";
       when X"09E" => sine <= X"000005FE";
       when X"09F" => sine <= X"000005BB";
       when X"0A0" => sine <= X"00000578";
       when X"0A1" => sine <= X"00000535";
       when X"0A2" => sine <= X"000004F1";
       when X"0A3" => sine <= X"000004AD";
       when X"0A4" => sine <= X"00000469";
       when X"0A5" => sine <= X"00000424";
       when X"0A6" => sine <= X"000003DE";
       when X"0A7" => sine <= X"00000399";
       when X"0A8" => sine <= X"00000353";
       when X"0A9" => sine <= X"0000030D";
       when X"0AA" => sine <= X"000002C7";
       when X"0AB" => sine <= X"00000280";
       when X"0AC" => sine <= X"0000023A";
       when X"0AD" => sine <= X"000001F3";
       when X"0AE" => sine <= X"000001AC";
       when X"0AF" => sine <= X"00000164";
       when X"0B0" => sine <= X"0000011D";
       when X"0B1" => sine <= X"000000D6";
       when X"0B2" => sine <= X"0000008E";
       when X"0B3" => sine <= X"00000047";
       when X"0B4" => sine <= X"00000000";
       when X"0B5" => sine <= X"FFFFFFB9";
       when X"0B6" => sine <= X"FFFFFF72";
       when X"0B7" => sine <= X"FFFFFF2A";
       when X"0B8" => sine <= X"FFFFFEE3";
       when X"0B9" => sine <= X"FFFFFE9C";
       when X"0BA" => sine <= X"FFFFFE54";
       when X"0BB" => sine <= X"FFFFFE0D";
       when X"0BC" => sine <= X"FFFFFDC6";
       when X"0BD" => sine <= X"FFFFFD80";
       when X"0BE" => sine <= X"FFFFFD39";
       when X"0BF" => sine <= X"FFFFFCF3";
       when X"0C0" => sine <= X"FFFFFCAD";
       when X"0C1" => sine <= X"FFFFFC67";
       when X"0C2" => sine <= X"FFFFFC22";
       when X"0C3" => sine <= X"FFFFFBDC";
       when X"0C4" => sine <= X"FFFFFB97";
       when X"0C5" => sine <= X"FFFFFB53";
       when X"0C6" => sine <= X"FFFFFB0F";
       when X"0C7" => sine <= X"FFFFFACB";
       when X"0C8" => sine <= X"FFFFFA88";
       when X"0C9" => sine <= X"FFFFFA45";
       when X"0CA" => sine <= X"FFFFFA02";
       when X"0CB" => sine <= X"FFFFF9C0";
       when X"0CC" => sine <= X"FFFFF97F";
       when X"0CD" => sine <= X"FFFFF93D";
       when X"0CE" => sine <= X"FFFFF8FD";
       when X"0CF" => sine <= X"FFFFF8BD";
       when X"0D0" => sine <= X"FFFFF87E";
       when X"0D1" => sine <= X"FFFFF83F";
       when X"0D2" => sine <= X"FFFFF800";
       when X"0D3" => sine <= X"FFFFF7C3";
       when X"0D4" => sine <= X"FFFFF786";
       when X"0D5" => sine <= X"FFFFF74A";
       when X"0D6" => sine <= X"FFFFF70E";
       when X"0D7" => sine <= X"FFFFF6D3";
       when X"0D8" => sine <= X"FFFFF699";
       when X"0D9" => sine <= X"FFFFF65F";
       when X"0DA" => sine <= X"FFFFF627";
       when X"0DB" => sine <= X"FFFFF5EF";
       when X"0DC" => sine <= X"FFFFF5B8";
       when X"0DD" => sine <= X"FFFFF581";
       when X"0DE" => sine <= X"FFFFF54C";
       when X"0DF" => sine <= X"FFFFF517";
       when X"0E0" => sine <= X"FFFFF4E3";
       when X"0E1" => sine <= X"FFFFF4B0";
       when X"0E2" => sine <= X"FFFFF47E";
       when X"0E3" => sine <= X"FFFFF44D";
       when X"0E4" => sine <= X"FFFFF41D";
       when X"0E5" => sine <= X"FFFFF3ED";
       when X"0E6" => sine <= X"FFFFF3BF";
       when X"0E7" => sine <= X"FFFFF391";
       when X"0E8" => sine <= X"FFFFF365";
       when X"0E9" => sine <= X"FFFFF339";
       when X"0EA" => sine <= X"FFFFF30F";
       when X"0EB" => sine <= X"FFFFF2E5";
       when X"0EC" => sine <= X"FFFFF2BD";
       when X"0ED" => sine <= X"FFFFF295";
       when X"0EE" => sine <= X"FFFFF26F";
       when X"0EF" => sine <= X"FFFFF24A";
       when X"0F0" => sine <= X"FFFFF225";
       when X"0F1" => sine <= X"FFFFF202";
       when X"0F2" => sine <= X"FFFFF1E0";
       when X"0F3" => sine <= X"FFFFF1BF";
       when X"0F4" => sine <= X"FFFFF19F";
       when X"0F5" => sine <= X"FFFFF180";
       when X"0F6" => sine <= X"FFFFF163";
       when X"0F7" => sine <= X"FFFFF146";
       when X"0F8" => sine <= X"FFFFF12B";
       when X"0F9" => sine <= X"FFFFF111";
       when X"0FA" => sine <= X"FFFFF0F8";
       when X"0FB" => sine <= X"FFFFF0E0";
       when X"0FC" => sine <= X"FFFFF0C9";
       when X"0FD" => sine <= X"FFFFF0B3";
       when X"0FE" => sine <= X"FFFFF09F";
       when X"0FF" => sine <= X"FFFFF08C";
       when X"100" => sine <= X"FFFFF07A";
       when X"101" => sine <= X"FFFFF069";
       when X"102" => sine <= X"FFFFF05A";
       when X"103" => sine <= X"FFFFF04C";
       when X"104" => sine <= X"FFFFF03F";
       when X"105" => sine <= X"FFFFF033";
       when X"106" => sine <= X"FFFFF028";
       when X"107" => sine <= X"FFFFF01F";
       when X"108" => sine <= X"FFFFF017";
       when X"109" => sine <= X"FFFFF010";
       when X"10A" => sine <= X"FFFFF00A";
       when X"10B" => sine <= X"FFFFF006";
       when X"10C" => sine <= X"FFFFF003";
       when X"10D" => sine <= X"FFFFF001";
       when X"10E" => sine <= X"FFFFF000";
       when X"10F" => sine <= X"FFFFF001";
       when X"110" => sine <= X"FFFFF003";
       when X"111" => sine <= X"FFFFF006";
       when X"112" => sine <= X"FFFFF00A";
       when X"113" => sine <= X"FFFFF010";
       when X"114" => sine <= X"FFFFF017";
       when X"115" => sine <= X"FFFFF01F";
       when X"116" => sine <= X"FFFFF028";
       when X"117" => sine <= X"FFFFF033";
       when X"118" => sine <= X"FFFFF03F";
       when X"119" => sine <= X"FFFFF04C";
       when X"11A" => sine <= X"FFFFF05A";
       when X"11B" => sine <= X"FFFFF069";
       when X"11C" => sine <= X"FFFFF07A";
       when X"11D" => sine <= X"FFFFF08C";
       when X"11E" => sine <= X"FFFFF09F";
       when X"11F" => sine <= X"FFFFF0B3";
       when X"120" => sine <= X"FFFFF0C9";
       when X"121" => sine <= X"FFFFF0E0";
       when X"122" => sine <= X"FFFFF0F8";
       when X"123" => sine <= X"FFFFF111";
       when X"124" => sine <= X"FFFFF12B";
       when X"125" => sine <= X"FFFFF146";
       when X"126" => sine <= X"FFFFF163";
       when X"127" => sine <= X"FFFFF180";
       when X"128" => sine <= X"FFFFF19F";
       when X"129" => sine <= X"FFFFF1BF";
       when X"12A" => sine <= X"FFFFF1E0";
       when X"12B" => sine <= X"FFFFF202";
       when X"12C" => sine <= X"FFFFF225";
       when X"12D" => sine <= X"FFFFF24A";
       when X"12E" => sine <= X"FFFFF26F";
       when X"12F" => sine <= X"FFFFF295";
       when X"130" => sine <= X"FFFFF2BD";
       when X"131" => sine <= X"FFFFF2E5";
       when X"132" => sine <= X"FFFFF30F";
       when X"133" => sine <= X"FFFFF339";
       when X"134" => sine <= X"FFFFF365";
       when X"135" => sine <= X"FFFFF391";
       when X"136" => sine <= X"FFFFF3BF";
       when X"137" => sine <= X"FFFFF3ED";
       when X"138" => sine <= X"FFFFF41D";
       when X"139" => sine <= X"FFFFF44D";
       when X"13A" => sine <= X"FFFFF47E";
       when X"13B" => sine <= X"FFFFF4B0";
       when X"13C" => sine <= X"FFFFF4E3";
       when X"13D" => sine <= X"FFFFF517";
       when X"13E" => sine <= X"FFFFF54C";
       when X"13F" => sine <= X"FFFFF581";
       when X"140" => sine <= X"FFFFF5B8";
       when X"141" => sine <= X"FFFFF5EF";
       when X"142" => sine <= X"FFFFF627";
       when X"143" => sine <= X"FFFFF65F";
       when X"144" => sine <= X"FFFFF699";
       when X"145" => sine <= X"FFFFF6D3";
       when X"146" => sine <= X"FFFFF70E";
       when X"147" => sine <= X"FFFFF74A";
       when X"148" => sine <= X"FFFFF786";
       when X"149" => sine <= X"FFFFF7C3";
       when X"14A" => sine <= X"FFFFF800";
       when X"14B" => sine <= X"FFFFF83F";
       when X"14C" => sine <= X"FFFFF87E";
       when X"14D" => sine <= X"FFFFF8BD";
       when X"14E" => sine <= X"FFFFF8FD";
       when X"14F" => sine <= X"FFFFF93D";
       when X"150" => sine <= X"FFFFF97F";
       when X"151" => sine <= X"FFFFF9C0";
       when X"152" => sine <= X"FFFFFA02";
       when X"153" => sine <= X"FFFFFA45";
       when X"154" => sine <= X"FFFFFA88";
       when X"155" => sine <= X"FFFFFACB";
       when X"156" => sine <= X"FFFFFB0F";
       when X"157" => sine <= X"FFFFFB53";
       when X"158" => sine <= X"FFFFFB97";
       when X"159" => sine <= X"FFFFFBDC";
       when X"15A" => sine <= X"FFFFFC22";
       when X"15B" => sine <= X"FFFFFC67";
       when X"15C" => sine <= X"FFFFFCAD";
       when X"15D" => sine <= X"FFFFFCF3";
       when X"15E" => sine <= X"FFFFFD39";
       when X"15F" => sine <= X"FFFFFD80";
       when X"160" => sine <= X"FFFFFDC6";
       when X"161" => sine <= X"FFFFFE0D";
       when X"162" => sine <= X"FFFFFE54";
       when X"163" => sine <= X"FFFFFE9C";
       when X"164" => sine <= X"FFFFFEE3";
       when X"165" => sine <= X"FFFFFF2A";
       when X"166" => sine <= X"FFFFFF72";
       when X"167" => sine <= X"FFFFFFB9";
       when X"168" => sine <= X"00000000";
       when others => sine <= X"FFFFFFFF";
       end case;
		 end if;
end process;
end Behavioral;